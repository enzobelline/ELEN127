module client()


